library ieee;
use ieee.std_logic_1164.all;

package Types is
    type std_logic_array is array (integer range <>) of std_logic_vector;
end package; -- Types
